// DDR3 Project Configuration Header File
`ifndef DDR3_DEFINES_VH
`define DDR3_DEFINES_VH

// 全局开关
`define SIMULATION
// `define DEBUG
// `define ONLINE

`endif  // DDR3_DEFINES_VH
