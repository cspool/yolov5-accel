// DDR3 Project Configuration Header File
`ifndef DDR3_DEFINES_VH
`define DDR3_DEFINES_VH

// `define SIMULATION
// `define CMD_DATA_SYNC
//`define DEBUG
`define ONLINE

`endif  // DDR3_DEFINES_VH
