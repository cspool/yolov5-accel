module product_add_bias_vecOp (
    clk,
    en,
    reset,
    mode,
    sum_mult_E_vector,  // pox res per channel
    bias_set,
    product_add_bias_vector  // pox res per channel
);

  parameter row_num_in_sa = 16;
  parameter column_num_in_sa = 16;
  parameter headroom = 8;
  parameter pixel_width_88 = 16 + headroom;
  parameter pixel_width_18 = 8 + headroom;
  parameter pe_parallel_pixel_88 = 2;
  parameter pe_parallel_weight_88 = 1;
  parameter pe_parallel_pixel_18 = 2;
  parameter pe_parallel_weight_18 = 2;
  parameter sa_row_num = 4;  //how many rows in conv core
  parameter sa_column_num = 3;  //how many columns in conv core
  parameter bias_width = 8;  //8 bit bias
  parameter bias_set_width = bias_width * pe_parallel_weight_18;  //16 bit
  parameter mult_P_width = 40;
  parameter sum_mult_E_vector_in_mult_P_width_width = mult_P_width * pe_parallel_weight_18 * pe_parallel_pixel_18 * column_num_in_sa;
  //40 bit * 32 pixels * 2 channel > 32 bit * 32 pixels * 2 channel > 40 bit * 32 pixels * 1 channel
  parameter sum_mult_E_vector_in_mult_P_width_width_88 = mult_P_width * pe_parallel_weight_88 * pe_parallel_pixel_88 * column_num_in_sa;
  parameter sum_mult_E_vector_in_mult_P_width_width_18_2 = mult_P_width * 1 * pe_parallel_pixel_18 * column_num_in_sa;
  parameter product_add_bias_vector_width = mult_P_width * pe_parallel_pixel_18 * pe_parallel_weight_18 * column_num_in_sa;
  parameter product_add_bias_vector_width_88 = mult_P_width * pe_parallel_pixel_88 * pe_parallel_weight_88 * column_num_in_sa;
  parameter product_add_bias_vector_width_18_2 = mult_P_width * pe_parallel_pixel_18 * 1 * column_num_in_sa;

  input clk, en, reset;
  input [3:0] mode;
  input [sum_mult_E_vector_in_mult_P_width_width - 1:0] sum_mult_E_vector;
  input [bias_set_width-1 : 0] bias_set;  //2 bias 16 bit, or 1 bias 8 bit
  output reg [product_add_bias_vector_width - 1:0] product_add_bias_vector;

  wire [bias_width-1 : 0] bias_88;
  wire [bias_width-1:0] bias_18_1, bias_18_2;

  wire [sum_mult_E_vector_in_mult_P_width_width_88 - 1 : 0] sum_mult_E_vector_88;
  wire [sum_mult_E_vector_in_mult_P_width_width_18_2 - 1 : 0] sum_mult_E_vector_18_1, sum_mult_E_vector_18_2;

  wire [product_add_bias_vector_width_88 - 1 : 0] product_add_bias_vector_88;
  wire [product_add_bias_vector_width_18_2 - 1 : 0] product_add_bias_vector_18_1, product_add_bias_vector_18_2;

  assign sum_mult_E_vector_88   = sum_mult_E_vector[sum_mult_E_vector_in_mult_P_width_width_88-1 : 0];
  assign sum_mult_E_vector_18_1 = sum_mult_E_vector[sum_mult_E_vector_in_mult_P_width_width_18_2-1 : 0];
  assign sum_mult_E_vector_18_2 = sum_mult_E_vector[sum_mult_E_vector_in_mult_P_width_width-1 : sum_mult_E_vector_in_mult_P_width_width_18_2];

  assign bias_88                = bias_set[bias_width-1 : 0];
  assign bias_18_1              = bias_88;
  assign bias_18_2              = bias_set[bias_set_width-1 : bias_width];

  genvar i;
  generate
    for (i = 0; i < pe_parallel_pixel_88 * pe_parallel_weight_88 * column_num_in_sa; i = i + 1) begin
      assign product_add_bias_vector_88[(i*mult_P_width)+:mult_P_width] =
          //sum * E
          sum_mult_E_vector_88[(i*mult_P_width)+:mult_P_width] +
          //bias
          {{(mult_P_width - bias_width) {bias_88[bias_width-1]}}, bias_88};  //bias_18_1 = bias_88
    end
    for (i = 0; i < pe_parallel_pixel_18 * 1 * column_num_in_sa; i = i + 1) begin
      assign product_add_bias_vector_18_1[(i*mult_P_width)+:mult_P_width] =
          //sum * E
          sum_mult_E_vector_18_1[(i*mult_P_width)+:mult_P_width] +
          //bias
          {{(mult_P_width - bias_width) {bias_18_1[bias_width-1]}}, bias_18_1};
    end
    for (i = 0; i < pe_parallel_pixel_18 * 1 * column_num_in_sa; i = i + 1) begin
      assign product_add_bias_vector_18_2[(i*mult_P_width)+:mult_P_width] =
          //sum * E
          sum_mult_E_vector_18_2[(i*mult_P_width)+:mult_P_width] +
          //bias
          {{(mult_P_width - bias_width) {bias_18_2[bias_width-1]}}, bias_18_2};
    end
  endgenerate

  always @(posedge clk) begin
    if (reset == 1'b1) begin
      product_add_bias_vector <= 0;
    end else if (en == 1'b1) begin
      product_add_bias_vector <=
      //mode 0
      (mode == 0) ? {{(product_add_bias_vector_width - product_add_bias_vector_width_88) {1'b0}}, product_add_bias_vector_88} :
      // mode 1
      (mode == 1) ? {product_add_bias_vector_18_2, product_add_bias_vector_18_1} : 0;
    end else begin
      product_add_bias_vector <= product_add_bias_vector;
    end
  end

endmodule
